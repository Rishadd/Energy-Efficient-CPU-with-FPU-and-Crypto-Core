
module mux_3_1(a,b,c,sel,y);

input [15:0] a,b,c;
input [1:0] sel ;
output [15:0] y ;
reg [15:0] mux_out ;

assign y = mux_out ;
always @(*)
    case(sel)
        2'b00 : mux_out=a ;
        2'b01 : mux_out=b ;
        2'b10 : mux_out=c ;
        default : mux_out=0;

    endcase
endmodule
